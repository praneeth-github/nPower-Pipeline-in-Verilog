module AND(
	input A,B,
	output O
	);
	
	assign O = A & B;

endmodule

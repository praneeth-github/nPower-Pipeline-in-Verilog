module OR(
	input A,B,
	output O
	);
	
	assign O = A | B;

endmodule
